
module BeagleGFPGABackend (
  input  clki
  );
endmodule
