module SegmentStepGenerator ();

endmodule
